`timescale 1ns/1ps
`include "assert.v"

module inst_br_test();
    reg     clk, rst;
    integer i  ;

    top top (clk,rst);

    always #1 clk = ~clk;
    initial begin
        $dumpfile("inst_br_test.vcd");
        $dumpvars;
        $dumpvars(0, top.openmips.regfile.regs[1]);
        $dumpvars(0, top.openmips.regfile.regs[3]);
        $dumpvars(0, top.openmips.regfile.regs[31]);

        $readmemh("../data/inst_br_test.txt", top.rom.memory, 0, 91);

        clk = 0;
        rst = 1;
        #20 rst = 0;
        #10 `AR(1,32'hxxxxxxxx);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'hxxxxxxxx);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000001);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000001);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000002);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000003);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000003);`AHI(32'h00000000);`ALO(32'h00000000);
        #2  `AR(1,32'h00000003);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000004);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000004);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000002C);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000005);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000005);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000006);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000007);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000008);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000008);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000009);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000A);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000A);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000002C);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000B);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000C);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000D);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000E);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000E);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000000F);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000010);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000010);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000011);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000012);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000013);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000013);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h0000014C);`AHI(32'h00000002);`ALO(32'h0000000E);
        #2  `AR(1,32'h00000014);`AHI(32'h00000002);`ALO(32'h0000000E);
        `PASS;
    end

endmodule